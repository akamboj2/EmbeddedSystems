
module pwm_system (
	clk_clk,
	pwm_0_conduit_end_export,
	reset_reset_n);	

	input		clk_clk;
	output		pwm_0_conduit_end_export;
	input		reset_reset_n;
endmodule
