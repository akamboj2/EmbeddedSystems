
module parport (
	clk_clk,
	parport_0_conduit_end_export,
	reset_reset_n);	

	input		clk_clk;
	inout	[7:0]	parport_0_conduit_end_export;
	input		reset_reset_n;
endmodule
